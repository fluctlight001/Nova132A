`include "lib/defines.vh"
module IC (
    input wire clk,
    input wire rst,
    input wire [`StallBus-1:0] stall
);
endmodule